context ieee_bit_context is
	library ieee;
	use ieee.numeric_bit.all;
end context ieee_bit_context;

context ieee_std_context is
	library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
end context ieee_std_context;